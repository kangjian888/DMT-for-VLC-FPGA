// =============================================================================
// Filename: LongTrainingSeqGen.v
// Author: 
// Email: jkangac@connect.ust.hk
// Affiliation: Hong Kong University of Science and Technology
// Description:
// -----------------------------------------------------------------------------
module LongTrainingSeqGen(
	input SYS_CLK,
	input PHY_RST,
	input LONG_ACK, //LONG training sequence sending enable
	output reg [27:0] LONG_TRAINING_SEQ,
	output reg [8:0] LONG_TRAINING_SEQ_INDEX,
	output reg LONG_TRAINING_SEQ_VALID
);

reg [1:0] frame_counter;
reg [7:0] symbol_counter;
reg [27:0] long_rom [127:0];

always @ (posedge SYS_CLK)
    begin
        if(PHY_RST)
        	begin
        		frame_counter <= 4'd0;
        		symbol_counter <= 5'd0;
        		LONG_TRAINING_SEQ <= 28'd0;
        		LONG_TRAINING_SEQ_VALID <= 1'b0;
        		LONG_TRAINING_SEQ_INDEX <= 9'd0;
        		long_rom[0] <=   28'b0000_0010_0100_0000_0000_0000_0000;
        		long_rom[1] <=   28'b0000_0010_0000_0011_1111_1011_1110;
        		long_rom[2] <=   28'b1111_1111_0110_1000_1110_1000_0110;
        		long_rom[3] <=   28'b0000_0000_1100_0111_1011_0010_1110;
        		long_rom[4] <=   28'b0000_0010_0100_1111_0110_1101_0010;
        		long_rom[5] <=   28'b1111_1110_1010_1011_1100_1100_0111;
        		long_rom[6] <=   28'b0000_0000_0100_0100_1001_1101_1101;
        		long_rom[7] <=   28'b0000_0001_1100_1000_1100_1001_0111;
        		long_rom[8] <=   28'b1111_1111_0001_0101_1000_0110_1110;
        		long_rom[9] <=   28'b0000_0000_0100_1101_0001_0011_1101;
        		long_rom[10] <=  28'b1111_1101_1100_1110_1000_0101_1000;
        		long_rom[11] <=  28'b1111_1111_0100_1011_0111_0101_0110;
        		long_rom[12] <=  28'b0000_0001_0111_1110_0011_1111_1111;
        		long_rom[13] <=  28'b0000_0001_1101_0100_1111_0101_1011;
        		long_rom[14] <=  28'b0000_0000_1010_1011_0111_0010_1110;
        		long_rom[15] <=  28'b0000_0000_1010_1111_0101_0000_1100;
        		long_rom[16] <=  28'b0000_0001_0100_0000_0000_0000_0000;
        		long_rom[17] <=  28'b1111_1110_1101_0111_0101_1000_1110;
        		long_rom[18] <=  28'b0000_0000_1110_0010_1011_0101_1000;
        		long_rom[19] <=  28'b1111_1110_1000_0000_1010_1010_0100;
        		long_rom[20] <=  28'b1111_1110_1000_1110_0001_1000_1000;
        		long_rom[21] <=  28'b1111_1110_0001_0101_0110_0010_1011;
        		long_rom[22] <=  28'b0000_0010_1100_0010_1100_1010_0100;
        		long_rom[23] <=  28'b1111_1111_0001_1110_0101_0100_1111;
        		long_rom[24] <=  28'b0000_0001_0100_0011_0111_1111_1110;
        		long_rom[25] <=  28'b1111_1111_0001_1101_1011_1010_0110;
        		long_rom[26] <=  28'b1111_1111_1100_1111_0001_1111_0011;
        		long_rom[27] <=  28'b0000_0010_0101_1100_0011_0011_0011;
        		long_rom[28] <=  28'b0000_0000_0100_0000_0101_0111_1000;
        		long_rom[29] <=  28'b1111_1101_1011_0010_0111_1001_0110;
        		long_rom[30] <=  28'b0000_0000_1000_1000_1111_1010_1101;
        		long_rom[31] <=  28'b1111_1111_1001_0001_1111_1000_0110;
        		long_rom[32] <=  28'b1111_1110_0100_0000_0000_0000_0000;
        		long_rom[33] <=  28'b1111_1110_0111_1110_1111_1111_1100;
        		long_rom[34] <=  28'b1111_1110_1001_1101_1101_1001_0100;
        		long_rom[35] <=  28'b0000_0001_0110_0001_0000_0101_1010;
        		long_rom[36] <=  28'b1111_1111_0110_0110_1010_0001_1100;
        		long_rom[37] <=  28'b0000_0000_0011_1110_1111_1000_0010;
        		long_rom[38] <=  28'b1111_1110_1001_0100_1110_1000_1110;
        		long_rom[39] <=  28'b1111_1101_1101_0111_0111_0011_0110;
        		long_rom[40] <=  28'b1111_1110_1010_0110_1000_1010_0001;
        		long_rom[41] <=  28'b0000_0000_1001_1011_1011_0000_0100;
        		long_rom[42] <=  28'b0000_0001_0101_0000_1101_0000_1101;
        		long_rom[43] <=  28'b1111_1111_1010_1011_1011_0010_1000;
        		long_rom[44] <=  28'b0000_0010_0010_1101_1111_1000_0110;
        		long_rom[45] <=  28'b1111_1111_1101_1001_0110_1100_0010;
        		long_rom[46] <=  28'b1111_1111_0000_1100_1100_0011_0001;
        		long_rom[47] <=  28'b0000_0010_0101_0101_0110_0101_0011;
        		long_rom[48] <=  28'b0000_0001_0100_0000_0000_0000_0000;
        		long_rom[49] <=  28'b0000_0001_0100_0010_1100_1011_0111;
        		long_rom[50] <=  28'b1111_1110_0001_0000_0010_0010_0100;
        		long_rom[51] <=  28'b0000_0001_0100_1101_0111_0011_1101;
        		long_rom[52] <=  28'b0000_0000_1100_0101_1010_1111_0010;
        		long_rom[53] <=  28'b1111_1110_1000_1111_1010_0110_1000;
        		long_rom[54] <=  28'b0000_0001_0010_0100_1101_1111_0011;
        		long_rom[55] <=  28'b1111_1110_1111_1001_1001_0110_0010;
        		long_rom[56] <=  28'b1111_1110_0000_0000_0110_1111_0100;
        		long_rom[57] <=  28'b1111_1110_1000_1111_0100_1100_0100;
        		long_rom[58] <=  28'b1111_1111_0010_0100_0110_1110_0011;
        		long_rom[59] <=  28'b0000_0001_1001_0100_1111_1001_0000;
        		long_rom[60] <=  28'b0000_0001_0000_1001_1001_1001_1010;
        		long_rom[61] <=  28'b0000_0000_0011_0000_0010_1100_0110;
        		long_rom[62] <=  28'b1111_1101_1111_0001_0010_0010_0000;
        		long_rom[63] <=  28'b0000_0000_0111_1110_0011_1111_0101;
        		long_rom[64] <=  28'b1111_1110_0100_0000_0000_0000_0000;
        		long_rom[65] <=  28'b0000_0000_0111_1110_0011_1111_0101;
        		long_rom[66] <=  28'b1111_1101_1111_0001_0010_0010_0000;
        		long_rom[67] <=  28'b0000_0000_0011_0000_0010_1100_0110;
        		long_rom[68] <=  28'b0000_0001_0000_1001_1001_1001_1010;
        		long_rom[69] <=  28'b0000_0001_1001_0100_1111_1001_0000;
        		long_rom[70] <=  28'b1111_1111_0010_0100_0110_1110_0011;
        		long_rom[71] <=  28'b1111_1110_1000_1111_0100_1100_0100;
        		long_rom[72] <=  28'b1111_1110_0000_0000_0110_1111_0100;
        		long_rom[73] <=  28'b1111_1110_1111_1001_1001_0110_0010;
        		long_rom[74] <=  28'b0000_0001_0010_0100_1101_1111_0011;
        		long_rom[75] <=  28'b1111_1110_1000_1111_1010_0110_1000;
        		long_rom[76] <=  28'b0000_0000_1100_0101_1010_1111_0010;
        		long_rom[77] <=  28'b0000_0001_0100_1101_0111_0011_1101;
        		long_rom[78] <=  28'b1111_1110_0001_0000_0010_0010_0100;
        		long_rom[79] <=  28'b0000_0001_0100_0010_1100_1011_0111;
        		long_rom[80] <=  28'b0000_0001_0100_0000_0000_0000_0000;
        		long_rom[81] <=  28'b0000_0010_0101_0101_0110_0101_0011;
        		long_rom[82] <=  28'b1111_1111_0000_1100_1100_0011_0001;
        		long_rom[83] <=  28'b1111_1111_1101_1001_0110_1100_0010;
        		long_rom[84] <=  28'b0000_0010_0010_1101_1111_1000_0110;
        		long_rom[85] <=  28'b1111_1111_1010_1011_1011_0010_1000;
        		long_rom[86] <=  28'b0000_0001_0101_0000_1101_0000_1101;
        		long_rom[87] <=  28'b0000_0000_1001_1011_1011_0000_0100;
        		long_rom[88] <=  28'b1111_1110_1010_0110_1000_1010_0001;
        		long_rom[89] <=  28'b1111_1101_1101_0111_0111_0011_0110;
        		long_rom[90] <=  28'b1111_1110_1001_0100_1110_1000_1110;
        		long_rom[91] <=  28'b0000_0000_0011_1110_1111_1000_0010;
        		long_rom[92] <=  28'b1111_1111_0110_0110_1010_0001_1100;
        		long_rom[93] <=  28'b0000_0001_0110_0001_0000_0101_1010;
        		long_rom[94] <=  28'b1111_1110_1001_1101_1101_1001_0100;
        		long_rom[95] <=  28'b1111_1110_0111_1110_1111_1111_1100;
        		long_rom[96] <=  28'b1111_1110_0100_0000_0000_0000_0000;
        		long_rom[97] <=  28'b1111_1111_1001_0001_1111_1000_0110;
        		long_rom[98] <=  28'b0000_0000_1000_1000_1111_1010_1101;
        		long_rom[99] <=  28'b1111_1101_1011_0010_0111_1001_0110;
        		long_rom[100] <= 28'b0000_0000_0100_0000_0101_0111_1000;
        		long_rom[101] <= 28'b0000_0010_0101_1100_0011_0011_0011;
        		long_rom[102] <= 28'b1111_1111_1100_1111_0001_1111_0011;
        		long_rom[103] <= 28'b1111_1111_0001_1101_1011_1010_0110;
        		long_rom[104] <= 28'b0000_0001_0100_0011_0111_1111_1110;
        		long_rom[105] <= 28'b1111_1111_0001_1110_0101_0100_1111;
        		long_rom[106] <= 28'b0000_0010_1100_0010_1100_1010_0100;
        		long_rom[107] <= 28'b1111_1110_0001_0101_0110_0010_1011;
        		long_rom[108] <= 28'b1111_1110_1000_1110_0001_1000_1000;
        		long_rom[109] <= 28'b1111_1110_1000_0000_1010_1010_0100;
        		long_rom[110] <= 28'b0000_0000_1110_0010_1011_0101_1000;
        		long_rom[111] <= 28'b1111_1110_1101_0111_0101_1000_1110;
        		long_rom[112] <= 28'b0000_0001_0100_0000_0000_0000_0000;
        		long_rom[113] <= 28'b0000_0000_1010_1111_0101_0000_1100;
        		long_rom[114] <= 28'b0000_0000_1010_1011_0111_0010_1110;
        		long_rom[115] <= 28'b0000_0001_1101_0100_1111_0101_1011;
        		long_rom[116] <= 28'b0000_0001_0111_1110_0011_1111_1111;
        		long_rom[117] <= 28'b1111_1111_0100_1011_0111_0101_0110;
        		long_rom[118] <= 28'b1111_1101_1100_1110_1000_0101_1000;
        		long_rom[119] <= 28'b0000_0000_0100_1101_0001_0011_1101;
        		long_rom[120] <= 28'b1111_1111_0001_0101_1000_0110_1110;
        		long_rom[121] <= 28'b0000_0001_1100_1000_1100_1001_0111;
        		long_rom[122] <= 28'b0000_0000_0100_0100_1001_1101_1101;
        		long_rom[123] <= 28'b1111_1110_1010_1011_1100_1100_0111;
        		long_rom[124] <= 28'b0000_0010_0100_1111_0110_1101_0010;
        		long_rom[125] <= 28'b0000_0000_1100_0111_1011_0010_1110;
        		long_rom[126] <= 28'b1111_1111_0110_1000_1110_1000_0110;
        		long_rom[127] <= 28'b0000_0010_0000_0011_1111_1011_1110;
        	end
        else
        	begin
        		if (LONG_ACK) 
        		    begin
        		    	if (frame_counter == 2'd0) 
        		    	    begin
        		    	    	if (symbol_counter == 8'd0) 
        		    	    	    begin
        		                        LONG_TRAINING_SEQ <= $signed(long_rom[symbol_counter+8'd96]) >>> 1;
        		                        LONG_TRAINING_SEQ_VALID <= 1'b1;
        		                        symbol_counter <= symbol_counter + 1'b1;
        		                        LONG_TRAINING_SEQ_INDEX <= LONG_TRAINING_SEQ_INDEX + 1'b1;          		    	    	        
        		    	    	    end
        		    	        else if (symbol_counter < 8'd31) 
        		    	            begin
        		                        LONG_TRAINING_SEQ <= long_rom[symbol_counter+8'd96];
        		                        LONG_TRAINING_SEQ_VALID <= 1'b1;
        		                        symbol_counter <= symbol_counter + 1'b1;
        		                        LONG_TRAINING_SEQ_INDEX <= LONG_TRAINING_SEQ_INDEX + 1'b1;        		    	                
        		    	            end
        		    	        else 
        		    	            begin
        		                        LONG_TRAINING_SEQ <= long_rom[symbol_counter+8'd96];
        		                        LONG_TRAINING_SEQ_VALID <= 1'b1;
        		                        symbol_counter <= 8'd0;
        		                        frame_counter <= frame_counter + 1'b1;
        		                        LONG_TRAINING_SEQ_INDEX <= LONG_TRAINING_SEQ_INDEX + 1'b1;        		    	                
        		    	            end
        		    	    end
        		        else if (frame_counter <= 2'd2) 
        		            begin
        		                if (symbol_counter < 8'd127) 
        		                    begin
        		                        LONG_TRAINING_SEQ <= long_rom[symbol_counter];
        		                        LONG_TRAINING_SEQ_VALID <= 1'b1;
        		                        symbol_counter <= symbol_counter + 1'b1;
        		                        LONG_TRAINING_SEQ_INDEX <= LONG_TRAINING_SEQ_INDEX + 1'b1;
        		                    end
        		                else 
        		                    begin
        		                        LONG_TRAINING_SEQ <= long_rom[symbol_counter];
        		                        LONG_TRAINING_SEQ_INDEX <= LONG_TRAINING_SEQ_INDEX + 1'b1;
        		                        LONG_TRAINING_SEQ_VALID <= 1'b1;
        		                        symbol_counter <= 8'd0;
        		                        frame_counter <= frame_counter + 1'b1;
        		                    end
        		            end
        		        else 
        		            begin
        		                frame_counter <= 4'd0;
        		                LONG_TRAINING_SEQ <= $signed(long_rom[symbol_counter]) >>> 1;
        		                LONG_TRAINING_SEQ_INDEX <= LONG_TRAINING_SEQ_INDEX + 1'b1;
        		            end
        		    end
        		else 
        		    begin
        		        LONG_TRAINING_SEQ <= 28'd0;
        		        LONG_TRAINING_SEQ_VALID <= 1'b0;
        		        LONG_TRAINING_SEQ_INDEX <= 9'd0;
        		        frame_counter <= 4'd0;
        		        symbol_counter <= 8'd0;
        		    end
        	end
    end

endmodule
